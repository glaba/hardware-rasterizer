module FinalProject();
	
	
	
endmodule