module UnitCircle(
	input logic clock,
	input logic[7:0] angle,
	output logic[17:0] x, y
);
	always_ff @ (posedge clock) begin 
		case (angle)
			8'd0: begin x <= 18'b000001000000000000; y <= 18'b000000000000000000; end
			8'd1: begin x <= 18'b000000111111111110; y <= 18'b000000000001101011; end
			8'd2: begin x <= 18'b000000111111111010; y <= 18'b000000000011010110; end
			8'd3: begin x <= 18'b000000111111110011; y <= 18'b000000000101000001; end
			8'd4: begin x <= 18'b000000111111101001; y <= 18'b000000000110101100; end
			8'd5: begin x <= 18'b000000111111011100; y <= 18'b000000001000010110; end
			8'd6: begin x <= 18'b000000111111001101; y <= 18'b000000001010000000; end
			8'd7: begin x <= 18'b000000111110111011; y <= 18'b000000001011101010; end
			8'd8: begin x <= 18'b000000111110100110; y <= 18'b000000001101010011; end
			8'd9: begin x <= 18'b000000111110001110; y <= 18'b000000001110111100; end
			8'd10: begin x <= 18'b000000111101110100; y <= 18'b000000010000100100; end
			8'd11: begin x <= 18'b000000111101010111; y <= 18'b000000010010001011; end
			8'd12: begin x <= 18'b000000111100110111; y <= 18'b000000010011110001; end
			8'd13: begin x <= 18'b000000111100010101; y <= 18'b000000010101010111; end
			8'd14: begin x <= 18'b000000111011101111; y <= 18'b000000010110111011; end
			8'd15: begin x <= 18'b000000111011001000; y <= 18'b000000011000011111; end
			8'd16: begin x <= 18'b000000111010011101; y <= 18'b000000011010000001; end
			8'd17: begin x <= 18'b000000111001110000; y <= 18'b000000011011100011; end
			8'd18: begin x <= 18'b000000111001000001; y <= 18'b000000011101000011; end
			8'd19: begin x <= 18'b000000111000001111; y <= 18'b000000011110100010; end
			8'd20: begin x <= 18'b000000110111011011; y <= 18'b000000011111111111; end
			8'd21: begin x <= 18'b000000110110100100; y <= 18'b000000100001011100; end
			8'd22: begin x <= 18'b000000110101101011; y <= 18'b000000100010110110; end
			8'd23: begin x <= 18'b000000110100101111; y <= 18'b000000100100001111; end
			8'd24: begin x <= 18'b000000110011110001; y <= 18'b000000100101100111; end
			8'd25: begin x <= 18'b000000110010110001; y <= 18'b000000100110111101; end
			8'd26: begin x <= 18'b000000110001101111; y <= 18'b000000101000010001; end
			8'd27: begin x <= 18'b000000110000101010; y <= 18'b000000101001100100; end
			8'd28: begin x <= 18'b000000101111100011; y <= 18'b000000101010110100; end
			8'd29: begin x <= 18'b000000101110011011; y <= 18'b000000101100000011; end
			8'd30: begin x <= 18'b000000101101010000; y <= 18'b000000101101010000; end
			8'd31: begin x <= 18'b000000101100000011; y <= 18'b000000101110011011; end
			8'd32: begin x <= 18'b000000101010110100; y <= 18'b000000101111100011; end
			8'd33: begin x <= 18'b000000101001100100; y <= 18'b000000110000101010; end
			8'd34: begin x <= 18'b000000101000010001; y <= 18'b000000110001101111; end
			8'd35: begin x <= 18'b000000100110111101; y <= 18'b000000110010110001; end
			8'd36: begin x <= 18'b000000100101100111; y <= 18'b000000110011110001; end
			8'd37: begin x <= 18'b000000100100001111; y <= 18'b000000110100101111; end
			8'd38: begin x <= 18'b000000100010110110; y <= 18'b000000110101101011; end
			8'd39: begin x <= 18'b000000100001011100; y <= 18'b000000110110100100; end
			8'd40: begin x <= 18'b000000100000000000; y <= 18'b000000110111011011; end
			8'd41: begin x <= 18'b000000011110100010; y <= 18'b000000111000001111; end
			8'd42: begin x <= 18'b000000011101000011; y <= 18'b000000111001000001; end
			8'd43: begin x <= 18'b000000011011100011; y <= 18'b000000111001110000; end
			8'd44: begin x <= 18'b000000011010000001; y <= 18'b000000111010011101; end
			8'd45: begin x <= 18'b000000011000011111; y <= 18'b000000111011001000; end
			8'd46: begin x <= 18'b000000010110111011; y <= 18'b000000111011101111; end
			8'd47: begin x <= 18'b000000010101010111; y <= 18'b000000111100010101; end
			8'd48: begin x <= 18'b000000010011110001; y <= 18'b000000111100110111; end
			8'd49: begin x <= 18'b000000010010001011; y <= 18'b000000111101010111; end
			8'd50: begin x <= 18'b000000010000100100; y <= 18'b000000111101110100; end
			8'd51: begin x <= 18'b000000001110111100; y <= 18'b000000111110001110; end
			8'd52: begin x <= 18'b000000001101010011; y <= 18'b000000111110100110; end
			8'd53: begin x <= 18'b000000001011101010; y <= 18'b000000111110111011; end
			8'd54: begin x <= 18'b000000001010000000; y <= 18'b000000111111001101; end
			8'd55: begin x <= 18'b000000001000010110; y <= 18'b000000111111011100; end
			8'd56: begin x <= 18'b000000000110101100; y <= 18'b000000111111101001; end
			8'd57: begin x <= 18'b000000000101000001; y <= 18'b000000111111110011; end
			8'd58: begin x <= 18'b000000000011010110; y <= 18'b000000111111111010; end
			8'd59: begin x <= 18'b000000000001101011; y <= 18'b000000111111111110; end
			8'd60: begin x <= 18'b000000000000000000; y <= 18'b000001000000000000; end
			8'd61: begin x <= 18'b111111111110010101; y <= 18'b000000111111111110; end
			8'd62: begin x <= 18'b111111111100101010; y <= 18'b000000111111111010; end
			8'd63: begin x <= 18'b111111111010111111; y <= 18'b000000111111110011; end
			8'd64: begin x <= 18'b111111111001010100; y <= 18'b000000111111101001; end
			8'd65: begin x <= 18'b111111110111101010; y <= 18'b000000111111011100; end
			8'd66: begin x <= 18'b111111110110000000; y <= 18'b000000111111001101; end
			8'd67: begin x <= 18'b111111110100010110; y <= 18'b000000111110111011; end
			8'd68: begin x <= 18'b111111110010101101; y <= 18'b000000111110100110; end
			8'd69: begin x <= 18'b111111110001000100; y <= 18'b000000111110001110; end
			8'd70: begin x <= 18'b111111101111011100; y <= 18'b000000111101110100; end
			8'd71: begin x <= 18'b111111101101110101; y <= 18'b000000111101010111; end
			8'd72: begin x <= 18'b111111101100001111; y <= 18'b000000111100110111; end
			8'd73: begin x <= 18'b111111101010101001; y <= 18'b000000111100010101; end
			8'd74: begin x <= 18'b111111101001000101; y <= 18'b000000111011101111; end
			8'd75: begin x <= 18'b111111100111100001; y <= 18'b000000111011001000; end
			8'd76: begin x <= 18'b111111100101111111; y <= 18'b000000111010011101; end
			8'd77: begin x <= 18'b111111100100011101; y <= 18'b000000111001110000; end
			8'd78: begin x <= 18'b111111100010111101; y <= 18'b000000111001000001; end
			8'd79: begin x <= 18'b111111100001011110; y <= 18'b000000111000001111; end
			8'd80: begin x <= 18'b111111100000000001; y <= 18'b000000110111011011; end
			8'd81: begin x <= 18'b111111011110100100; y <= 18'b000000110110100100; end
			8'd82: begin x <= 18'b111111011101001010; y <= 18'b000000110101101011; end
			8'd83: begin x <= 18'b111111011011110001; y <= 18'b000000110100101111; end
			8'd84: begin x <= 18'b111111011010011001; y <= 18'b000000110011110001; end
			8'd85: begin x <= 18'b111111011001000011; y <= 18'b000000110010110001; end
			8'd86: begin x <= 18'b111111010111101111; y <= 18'b000000110001101111; end
			8'd87: begin x <= 18'b111111010110011100; y <= 18'b000000110000101010; end
			8'd88: begin x <= 18'b111111010101001100; y <= 18'b000000101111100011; end
			8'd89: begin x <= 18'b111111010011111101; y <= 18'b000000101110011011; end
			8'd90: begin x <= 18'b111111010010110000; y <= 18'b000000101101010000; end
			8'd91: begin x <= 18'b111111010001100101; y <= 18'b000000101100000011; end
			8'd92: begin x <= 18'b111111010000011101; y <= 18'b000000101010110100; end
			8'd93: begin x <= 18'b111111001111010110; y <= 18'b000000101001100100; end
			8'd94: begin x <= 18'b111111001110010001; y <= 18'b000000101000010001; end
			8'd95: begin x <= 18'b111111001101001111; y <= 18'b000000100110111101; end
			8'd96: begin x <= 18'b111111001100001111; y <= 18'b000000100101100111; end
			8'd97: begin x <= 18'b111111001011010001; y <= 18'b000000100100001111; end
			8'd98: begin x <= 18'b111111001010010101; y <= 18'b000000100010110110; end
			8'd99: begin x <= 18'b111111001001011100; y <= 18'b000000100001011100; end
			8'd100: begin x <= 18'b111111001000100101; y <= 18'b000000011111111111; end
			8'd101: begin x <= 18'b111111000111110001; y <= 18'b000000011110100010; end
			8'd102: begin x <= 18'b111111000110111111; y <= 18'b000000011101000011; end
			8'd103: begin x <= 18'b111111000110010000; y <= 18'b000000011011100011; end
			8'd104: begin x <= 18'b111111000101100011; y <= 18'b000000011010000001; end
			8'd105: begin x <= 18'b111111000100111000; y <= 18'b000000011000011111; end
			8'd106: begin x <= 18'b111111000100010001; y <= 18'b000000010110111011; end
			8'd107: begin x <= 18'b111111000011101011; y <= 18'b000000010101010111; end
			8'd108: begin x <= 18'b111111000011001001; y <= 18'b000000010011110001; end
			8'd109: begin x <= 18'b111111000010101001; y <= 18'b000000010010001011; end
			8'd110: begin x <= 18'b111111000010001100; y <= 18'b000000010000100100; end
			8'd111: begin x <= 18'b111111000001110010; y <= 18'b000000001110111100; end
			8'd112: begin x <= 18'b111111000001011010; y <= 18'b000000001101010011; end
			8'd113: begin x <= 18'b111111000001000101; y <= 18'b000000001011101010; end
			8'd114: begin x <= 18'b111111000000110011; y <= 18'b000000001010000000; end
			8'd115: begin x <= 18'b111111000000100100; y <= 18'b000000001000010110; end
			8'd116: begin x <= 18'b111111000000010111; y <= 18'b000000000110101100; end
			8'd117: begin x <= 18'b111111000000001101; y <= 18'b000000000101000001; end
			8'd118: begin x <= 18'b111111000000000110; y <= 18'b000000000011010110; end
			8'd119: begin x <= 18'b111111000000000010; y <= 18'b000000000001101011; end
			8'd120: begin x <= 18'b111111000000000000; y <= 18'b000000000000000000; end
			8'd121: begin x <= 18'b111111000000000010; y <= 18'b111111111110010101; end
			8'd122: begin x <= 18'b111111000000000110; y <= 18'b111111111100101010; end
			8'd123: begin x <= 18'b111111000000001101; y <= 18'b111111111010111111; end
			8'd124: begin x <= 18'b111111000000010111; y <= 18'b111111111001010100; end
			8'd125: begin x <= 18'b111111000000100100; y <= 18'b111111110111101010; end
			8'd126: begin x <= 18'b111111000000110011; y <= 18'b111111110110000000; end
			8'd127: begin x <= 18'b111111000001000101; y <= 18'b111111110100010110; end
			8'd128: begin x <= 18'b111111000001011010; y <= 18'b111111110010101101; end
			8'd129: begin x <= 18'b111111000001110010; y <= 18'b111111110001000100; end
			8'd130: begin x <= 18'b111111000010001100; y <= 18'b111111101111011100; end
			8'd131: begin x <= 18'b111111000010101001; y <= 18'b111111101101110101; end
			8'd132: begin x <= 18'b111111000011001001; y <= 18'b111111101100001111; end
			8'd133: begin x <= 18'b111111000011101011; y <= 18'b111111101010101001; end
			8'd134: begin x <= 18'b111111000100010001; y <= 18'b111111101001000101; end
			8'd135: begin x <= 18'b111111000100111000; y <= 18'b111111100111100001; end
			8'd136: begin x <= 18'b111111000101100011; y <= 18'b111111100101111111; end
			8'd137: begin x <= 18'b111111000110010000; y <= 18'b111111100100011101; end
			8'd138: begin x <= 18'b111111000110111111; y <= 18'b111111100010111101; end
			8'd139: begin x <= 18'b111111000111110001; y <= 18'b111111100001011110; end
			8'd140: begin x <= 18'b111111001000100101; y <= 18'b111111100000000000; end
			8'd141: begin x <= 18'b111111001001011100; y <= 18'b111111011110100100; end
			8'd142: begin x <= 18'b111111001010010101; y <= 18'b111111011101001010; end
			8'd143: begin x <= 18'b111111001011010001; y <= 18'b111111011011110001; end
			8'd144: begin x <= 18'b111111001100001111; y <= 18'b111111011010011001; end
			8'd145: begin x <= 18'b111111001101001111; y <= 18'b111111011001000011; end
			8'd146: begin x <= 18'b111111001110010001; y <= 18'b111111010111101111; end
			8'd147: begin x <= 18'b111111001111010110; y <= 18'b111111010110011100; end
			8'd148: begin x <= 18'b111111010000011101; y <= 18'b111111010101001100; end
			8'd149: begin x <= 18'b111111010001100101; y <= 18'b111111010011111101; end
			8'd150: begin x <= 18'b111111010010110000; y <= 18'b111111010010110000; end
			8'd151: begin x <= 18'b111111010011111101; y <= 18'b111111010001100101; end
			8'd152: begin x <= 18'b111111010101001100; y <= 18'b111111010000011101; end
			8'd153: begin x <= 18'b111111010110011100; y <= 18'b111111001111010110; end
			8'd154: begin x <= 18'b111111010111101111; y <= 18'b111111001110010001; end
			8'd155: begin x <= 18'b111111011001000011; y <= 18'b111111001101001111; end
			8'd156: begin x <= 18'b111111011010011001; y <= 18'b111111001100001111; end
			8'd157: begin x <= 18'b111111011011110001; y <= 18'b111111001011010001; end
			8'd158: begin x <= 18'b111111011101001010; y <= 18'b111111001010010101; end
			8'd159: begin x <= 18'b111111011110100100; y <= 18'b111111001001011100; end
			8'd160: begin x <= 18'b111111100000000000; y <= 18'b111111001000100101; end
			8'd161: begin x <= 18'b111111100001011110; y <= 18'b111111000111110001; end
			8'd162: begin x <= 18'b111111100010111101; y <= 18'b111111000110111111; end
			8'd163: begin x <= 18'b111111100100011101; y <= 18'b111111000110010000; end
			8'd164: begin x <= 18'b111111100101111111; y <= 18'b111111000101100011; end
			8'd165: begin x <= 18'b111111100111100001; y <= 18'b111111000100111000; end
			8'd166: begin x <= 18'b111111101001000101; y <= 18'b111111000100010001; end
			8'd167: begin x <= 18'b111111101010101001; y <= 18'b111111000011101011; end
			8'd168: begin x <= 18'b111111101100001111; y <= 18'b111111000011001001; end
			8'd169: begin x <= 18'b111111101101110101; y <= 18'b111111000010101001; end
			8'd170: begin x <= 18'b111111101111011100; y <= 18'b111111000010001100; end
			8'd171: begin x <= 18'b111111110001000100; y <= 18'b111111000001110010; end
			8'd172: begin x <= 18'b111111110010101101; y <= 18'b111111000001011010; end
			8'd173: begin x <= 18'b111111110100010110; y <= 18'b111111000001000101; end
			8'd174: begin x <= 18'b111111110110000000; y <= 18'b111111000000110011; end
			8'd175: begin x <= 18'b111111110111101010; y <= 18'b111111000000100100; end
			8'd176: begin x <= 18'b111111111001010100; y <= 18'b111111000000010111; end
			8'd177: begin x <= 18'b111111111010111111; y <= 18'b111111000000001101; end
			8'd178: begin x <= 18'b111111111100101010; y <= 18'b111111000000000110; end
			8'd179: begin x <= 18'b111111111110010101; y <= 18'b111111000000000010; end
			8'd180: begin x <= 18'b000000000000000000; y <= 18'b111111000000000000; end
			8'd181: begin x <= 18'b000000000001101011; y <= 18'b111111000000000010; end
			8'd182: begin x <= 18'b000000000011010110; y <= 18'b111111000000000110; end
			8'd183: begin x <= 18'b000000000101000001; y <= 18'b111111000000001101; end
			8'd184: begin x <= 18'b000000000110101100; y <= 18'b111111000000010111; end
			8'd185: begin x <= 18'b000000001000010110; y <= 18'b111111000000100100; end
			8'd186: begin x <= 18'b000000001010000000; y <= 18'b111111000000110011; end
			8'd187: begin x <= 18'b000000001011101010; y <= 18'b111111000001000101; end
			8'd188: begin x <= 18'b000000001101010011; y <= 18'b111111000001011010; end
			8'd189: begin x <= 18'b000000001110111100; y <= 18'b111111000001110010; end
			8'd190: begin x <= 18'b000000010000100100; y <= 18'b111111000010001100; end
			8'd191: begin x <= 18'b000000010010001011; y <= 18'b111111000010101001; end
			8'd192: begin x <= 18'b000000010011110001; y <= 18'b111111000011001001; end
			8'd193: begin x <= 18'b000000010101010111; y <= 18'b111111000011101011; end
			8'd194: begin x <= 18'b000000010110111011; y <= 18'b111111000100010001; end
			8'd195: begin x <= 18'b000000011000011111; y <= 18'b111111000100111000; end
			8'd196: begin x <= 18'b000000011010000001; y <= 18'b111111000101100011; end
			8'd197: begin x <= 18'b000000011011100011; y <= 18'b111111000110010000; end
			8'd198: begin x <= 18'b000000011101000011; y <= 18'b111111000110111111; end
			8'd199: begin x <= 18'b000000011110100010; y <= 18'b111111000111110001; end
			8'd200: begin x <= 18'b000000100000000000; y <= 18'b111111001000100101; end
			8'd201: begin x <= 18'b000000100001011100; y <= 18'b111111001001011100; end
			8'd202: begin x <= 18'b000000100010110110; y <= 18'b111111001010010101; end
			8'd203: begin x <= 18'b000000100100001111; y <= 18'b111111001011010001; end
			8'd204: begin x <= 18'b000000100101100111; y <= 18'b111111001100001111; end
			8'd205: begin x <= 18'b000000100110111101; y <= 18'b111111001101001111; end
			8'd206: begin x <= 18'b000000101000010001; y <= 18'b111111001110010001; end
			8'd207: begin x <= 18'b000000101001100100; y <= 18'b111111001111010110; end
			8'd208: begin x <= 18'b000000101010110100; y <= 18'b111111010000011101; end
			8'd209: begin x <= 18'b000000101100000011; y <= 18'b111111010001100101; end
			8'd210: begin x <= 18'b000000101101010000; y <= 18'b111111010010110000; end
			8'd211: begin x <= 18'b000000101110011011; y <= 18'b111111010011111101; end
			8'd212: begin x <= 18'b000000101111100011; y <= 18'b111111010101001100; end
			8'd213: begin x <= 18'b000000110000101010; y <= 18'b111111010110011100; end
			8'd214: begin x <= 18'b000000110001101111; y <= 18'b111111010111101111; end
			8'd215: begin x <= 18'b000000110010110001; y <= 18'b111111011001000011; end
			8'd216: begin x <= 18'b000000110011110001; y <= 18'b111111011010011001; end
			8'd217: begin x <= 18'b000000110100101111; y <= 18'b111111011011110001; end
			8'd218: begin x <= 18'b000000110101101011; y <= 18'b111111011101001010; end
			8'd219: begin x <= 18'b000000110110100100; y <= 18'b111111011110100100; end
			8'd220: begin x <= 18'b000000110111011011; y <= 18'b111111100000000000; end
			8'd221: begin x <= 18'b000000111000001111; y <= 18'b111111100001011110; end
			8'd222: begin x <= 18'b000000111001000001; y <= 18'b111111100010111101; end
			8'd223: begin x <= 18'b000000111001110000; y <= 18'b111111100100011101; end
			8'd224: begin x <= 18'b000000111010011101; y <= 18'b111111100101111111; end
			8'd225: begin x <= 18'b000000111011001000; y <= 18'b111111100111100001; end
			8'd226: begin x <= 18'b000000111011101111; y <= 18'b111111101001000101; end
			8'd227: begin x <= 18'b000000111100010101; y <= 18'b111111101010101001; end
			8'd228: begin x <= 18'b000000111100110111; y <= 18'b111111101100001111; end
			8'd229: begin x <= 18'b000000111101010111; y <= 18'b111111101101110101; end
			8'd230: begin x <= 18'b000000111101110100; y <= 18'b111111101111011100; end
			8'd231: begin x <= 18'b000000111110001110; y <= 18'b111111110001000100; end
			8'd232: begin x <= 18'b000000111110100110; y <= 18'b111111110010101101; end
			8'd233: begin x <= 18'b000000111110111011; y <= 18'b111111110100010110; end
			8'd234: begin x <= 18'b000000111111001101; y <= 18'b111111110110000000; end
			8'd235: begin x <= 18'b000000111111011100; y <= 18'b111111110111101010; end
			8'd236: begin x <= 18'b000000111111101001; y <= 18'b111111111001010100; end
			8'd237: begin x <= 18'b000000111111110011; y <= 18'b111111111010111111; end
			8'd238: begin x <= 18'b000000111111111010; y <= 18'b111111111100101010; end
			8'd239: begin x <= 18'b000000111111111110; y <= 18'b111111111110010101; end
		endcase 
	end 

endmodule 

module Motion(
	input logic clock, reset, update_position,
	input logic move_left, move_right, move_up, move_down, 
	input logic turn_left, turn_right, turn_up, turn_down,
	input logic move_forward, move_backward,
	output logic[17:0] camera_origin[2:0], u_vec[2:0], v_vec[2:0], n_vec[2:0], light_vec[2:0]
);
	logic[7:0] angle, angle_in;
	logic[17:0] x, y;
	logic[3:0] update_angle; // To prevent the angle from changing too fast
	UnitCircle uc(.clock, .angle, .x, .y);

	logic[17:0] u_displacement[2:0], v_displacement[2:0], n_displacement[2:0], displacement[2:0];
	always_ff @ (posedge clock) begin 
		u_vec[2] <= x; u_vec[1] <= 18'd0; u_vec[0] <= y;
		n_vec[2] <= ~y + 18'd1; n_vec[1] <= 18'd0; n_vec[0] <= x;
		// It's like you're shining a flashlight
		light_vec[2] <= ~y + 18'd1; light_vec[1] <= 18'd0; light_vec[0] <= x;
		
		if (reset) begin 
			angle <= 8'd0;	
			update_angle <= 4'd0;

			// (0, 0, -1)
			v_vec[2] <= 18'd0; v_vec[1] <= {6'd1, 12'd0}; v_vec[0] <= 18'd0;

			// (0, 0, -10)
			camera_origin[2] <= 18'd0; camera_origin[1] <= 18'd0; camera_origin[0] <= {6'b110110, 12'd0};
		end 
		else begin 
			if (update_position & (update_angle == 4'd0)) angle <= angle_in;
			else                                          angle <= angle;

			if (update_angle == 4'd9) update_angle <= 4'd0;
			else                      update_angle <= update_angle + 4'd1;

			for (int i = 0; i < 3; i++) begin 
				v_vec[i] <= v_vec[i];

				if (update_position) begin 
					camera_origin[i] <= camera_origin[i] + displacement[i];
				end 
				else begin 
					camera_origin[i] <= camera_origin[i];
				end 
			end 
		end 
	end 

	always_comb begin 
		if (turn_right) begin 
			if (angle == 8'd0) angle_in = 8'd239;
			else               angle_in = angle - 8'd1;
		end 
		else if (turn_left) begin 
			if (angle == 8'd239) angle_in = 8'd0;
			else                 angle_in = angle + 8'd1;
		end 
		else begin 
			angle_in = angle;
		end 

		for (int i = 0; i < 3; i++) begin 
			if (move_left)       u_displacement[i] = ~{{6{u_vec[i][17]}}, u_vec[i][17:6]} + 18'd1;
			else if (move_right) u_displacement[i] = {{6{u_vec[i][17]}}, u_vec[i][17:6]};
			else                 u_displacement[i] = 18'd0;

			if (move_up)        v_displacement[i] = ~{{6{v_vec[i][17]}}, v_vec[i][17:6]} + 18'd1;
			else if (move_down) v_displacement[i] = {{6{v_vec[i][17]}}, v_vec[i][17:6]};
			else                v_displacement[i] = 18'd0;

			if (move_forward)       n_displacement[i] = {{6{n_vec[i][17]}}, n_vec[i][17:6]};
			else if (move_backward) n_displacement[i] = ~{{6{n_vec[i][17]}}, n_vec[i][17:6]} + 18'd1;
			else                    n_displacement[i] = 18'd0;

			displacement[i] = u_displacement[i] + v_displacement[i] + n_displacement[i];
		end 
	end 
endmodule 